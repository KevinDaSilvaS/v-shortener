module structs

pub enum FileFormats {
	html
	json
	text
}