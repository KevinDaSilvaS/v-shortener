module structs

pub struct CreatedLink {
    pub: link_name string
         creation_date string
}