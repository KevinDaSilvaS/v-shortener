module structs

pub type Response = CreatedLink | string | ApiError