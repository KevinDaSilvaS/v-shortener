module structs

pub struct ApiError {
	message string
}