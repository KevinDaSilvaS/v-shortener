module requests

pub struct CreateLinkRequest {
	pub: link_name string
}